library verilog;
use verilog.vl_types.all;
entity testing_counter_vlg_vec_tst is
end testing_counter_vlg_vec_tst;
